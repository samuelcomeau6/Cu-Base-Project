`timescale 1ns / 1ns
///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////
///
/// Top-Level Verilog Module
///
/// Only include pins the design is actually using.  Make sure that the pin is
/// given the correct direction: input vs. output vs. inout
///
///////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////
module Cu_tb (
);
    reg clk;
    reg rst_n;
    reg[7:0] leg;
    reg usb_rx;
    reg usb_tx;
    always #5 clk=~clk;
    initial begin
        #10000000
        $display("Test Sat");
        $finish;
    end
endmodule
